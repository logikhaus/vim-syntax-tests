/* Standard IEEE P1076.6 directives. */
/*rtl_synthesison*/			-- not marked up.
/*rtl_synthesisoff*/		-- not marked up.
/*rtl_synthesis on*/
/*rtl_synthesis off*/
/* RTL_SYNTHESIS ON */
/* RTL_SYNTHESIS OFF */
/* rtl_synthesis on */
/* rtl_synthesis off */
/* rtl_synthesis	on */
/* rtl_synthesis	off */
	/* rtl_synthesis on */
	/* rtl_synthesis off */
/*rtl_syn on*/
/*rtl_syn off*/
/* RTL_SYN ON */
/* RTL_SYN OFF */
/* rtl_syn on */
/* rtl_syn off */
/* rtl_syn	on */
/* rtl_syn	off */
	/* rtl_syn on */
	/* rtl_syn off */
--rtl_synthesison			-- not marked up.
--rtl_synthesisoff			-- not marked up.
--RTL_SYNTHESIS ON
--RTL_SYNTHESIS OFF
--rtl_synthesis on
--rtl_synthesis off
-- rtl_synthesis on
-- rtl_synthesis off
-- rtl_synthesis on 
-- rtl_synthesis off 
-- rtl_synthesis	on
-- rtl_synthesis	off
	-- rtl_synthesis on 
	-- rtl_synthesis off
--rtl_synon					-- not marked up.
--rtl_synoff				-- not marked up.
--RTL_SYN ON
--RTL_SYN OFF
--rtl_syn on
--rtl_syn off
-- rtl_syn on
-- rtl_syn off
-- rtl_syn on 
-- rtl_syn off 
-- rtl_syn	on
-- rtl_syn	off
	-- rtl_syn on 
	-- rtl_syn off

/* Industry-standard directives. */

/*synthesistranslate_on*/				-- not marked up.
/*synthesistranslate_off*/				-- not marked up.
/*synthesis translate_on*/
/*synthesis translate_off*/
/* synthesis translate_on */
/* synthesis translate_off */
/* synthesis	translate_on */
/* synthesis	translate_off */
	/* synthesis translate_on */
	/* synthesis translate_off */
--synthesistranslate_on					-- not marked up.
--synthesistranslate_off				-- not marked up.
--synthesis translate_on
--synthesis translate_off
-- synthesis translate_on
-- synthesis translate_off
-- synthesis translate_on 
-- synthesis translate_off 
-- synthesis	translate_on
-- synthesis	translate_off
	-- synthesis translate_on 
	-- synthesis translate_off

/*simulationtranslate_on*/				-- not marked up.
/*simulationtranslate_off*/				-- not marked up.
/*simulation translate_on*/
/*simulation translate_off*/
/* simulation translate_on */
/* simulation translate_off */
/* simulation	translate_on */
/* simulation	translate_off */
	/* simulation translate_on */
	/* simulation translate_off */
--simulationtranslate_on				-- not marked up.
--simulationtranslate_off				-- not marked up.
--simulation translate_on
--simulation translate_off
-- simulation translate_on
-- simulation translate_off
-- simulation translate_on 
-- simulation translate_off 
-- simulation	translate_on
-- simulation	translate_off
	-- simulation translate_on
	-- simulation translate_off

/*synopsystranslate_on*/				-- not marked up.
/*synopsystranslate_off*/				-- not marked up.
/*synopsys translate_on*/
/*synopsys translate_off*/
/* synopsys translate_on */
/* synopsys translate_off */
/* synopsys	translate_on */
/* synopsys	translate_off */
	/* synopsys translate_on */
	/* synopsys translate_off */
--synopsystranslate_on					-- not marked up.
--synopsystranslate_off					-- not marked up.
--synopsys translate_on
--synopsys translate_off
-- synopsys translate_on
-- synopsys translate_off
-- synopsys translate_on 
-- synopsys translate_off 
-- synopsys	translate_on
-- synopsys	translate_off
	-- synopsys translate_on
	-- synopsys translate_off

/*pragmatranslate_on*/					-- not marked up.
/*pragmatranslate_off*/					-- not marked up.
/*pragma translate_on*/
/*pragma translate_off*/
/* pragma translate_on */
/* pragma translate_off */
/* pragma	translate_on */
/* pragma	translate_off */
	/* pragma translate_on */
	/* pragma translate_off */
--pragmatranslate_on					-- not marked up.
--pragmatranslate_off					-- not marked up.
--pragma translate_on
--pragma translate_off
-- pragma translate_on
-- pragma translate_off
-- pragma translate_on 
-- pragma translate_off 
-- pragma	translate_on
-- pragma	translate_off
-- pragma translate_on
-- pragma translate_off
	-- pragma translate_on
	-- pragma translate_off

/*pragmasynthesis_on*/					-- not marked up.
/*pragmasynthesis_off*/					-- not marked up.
/*pragma synthesis_on*/
/*pragma synthesis_off*/
/* pragma synthesis_on */
/* pragma synthesis_off */
/* pragma	synthesis_on */
/* pragma	synthesis_off */
	/* pragma synthesis_on */
	/* pragma synthesis_off */
--pragmasynthesis_on					-- not marked up.
--pragmasynthesis_off					-- not marked up.
--pragma synthesis_on
--pragma synthesis_off
-- pragma synthesis_on
-- pragma synthesis_off
-- pragma synthesis_on 
-- pragma synthesis_off 
-- pragma	synthesis_on
-- pragma	synthesis_off
-- pragma synthesis_on
-- pragma synthesis_off
	-- pragma synthesis_on
	-- pragma synthesis_off
